���/      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��h2�f8�����R�(KhHNNNJ����J����K t�b�C              �?�t�bhLh&�scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hxhGK ��hyhGK��hzhGK��h{hXK��h|hXK ��h}hGK(��h~hXK0��uK8KKt�b�Bh                              @�\��N��?             C@������������������������       �                     1@       
                    �?���N8�?             5@                          �g@�����H�?             "@������������������������       �                     @                          �@@�q�q�?             @������������������������       �                     �?       	                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�t�b�values�h(h+K ��h-��R�(KKKK��hX�C�      2@      4@      1@              �?      4@      �?       @              @      �?       @              �?      �?      �?      �?                      �?              (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @�\��N��?             C@������������������������       �        
             *@                            @ �o_��?             9@                           @      �?             ,@                          �@@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      4@      2@      *@              @      2@      @      @      @       @      @                       @              @              &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @D�n�3�?             C@                          �d@�8��8��?             8@                          �d@����X�?             @                           N@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             1@������������������������       �        	             ,@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�      6@      0@      6@       @      @       @      @      �?      @                      �?              �?      1@                      ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                              @p�ݯ��?             C@������������������������       �                     $@       
                     @؇���X�?             <@       	                   �g@���|���?             &@                          �@@�<ݚ�?             "@                          �:@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     1@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      ,@      8@      $@              @      8@      @      @       @      @       @      @              @       @                      @       @                      1@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @      �?             C@������������������������       �        
             0@       
                   �g@��2(&�?             6@       	                   �@@�IєX�?             1@                         ��e@r�q��?             @������������������������       �                     @                         �5g@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@                            @���Q��?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      3@      3@      0@              @      3@      �?      0@      �?      @              @      �?       @      �?                       @              &@       @      @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                             6@      �?             C@������������������������       �                     @                           �?4���C�?            �@@������������������������       �                     "@                            @�q�q�?             8@������������������������       �                     @       
                   �@@�����?             5@       	                     @����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     ,@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      3@      3@      @              ,@      3@      "@              @      3@      @               @      3@       @      @       @                      @              ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                            �h@D�n�3�?             C@                            @�q�q�?            �@@                            @d}h���?             ,@������������������������       �                      @       
                   �g@      �?             @       	                  �%g@      �?             @                          �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             3@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      0@      6@      &@      6@      &@      @       @              @      @      �?      @      �?      �?      �?                      �?               @       @                      3@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�BH                              @D�n�3�?             C@������������������������       �                     "@                           C@>���Rp�?             =@                            @j���� �?             1@                          �g@�z�G��?             $@       	                    �?���Q��?             @                          �:@      �?              @������������������������       �                     �?������������������������       �                     �?
                         �%g@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      0@      6@      "@              @      6@      @      $@      @      @       @      @      �?      �?              �?      �?              �?       @      �?                       @      @                      @              (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                             6@�\��N��?             C@������������������������       �                     @                            @����e��?            �@@������������������������       �                     &@       
                     @�C��2(�?             6@                           �?�<ݚ�?             "@������������������������       �                     �?       	                   �@@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        	             *@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      2@      4@      @              *@      4@      &@               @      4@       @      @      �?              �?      @      �?                      @              *@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @p�ݯ��?             C@������������������������       �        
             3@                          �@@�d�����?             3@                            @X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      8@      ,@      3@              @      ,@      @      @      @                      @              $@�t�bubhhubehhub.